module AND_Gate(
  input A,
  input B,
  output Y);
  
  assign Y = A&&B; // Y is the opposite of A
  
endmodule
